module regfile(
    input clk,
    input reg_write,
    input [4:0] rs1,
    input [4:0] rs2,
    input [4:0] rd,
    input [31:0] wd,
    output [31:0] rd1,
    output [31:0] rd2
);

reg [31:0] regs [31:0];

// Read (combinational)
assign rd1 = (rs1 == 0) ? 32'b0 : regs[rs1];
assign rd2 = (rs2 == 0) ? 32'b0 : regs[rs2];

// Write (sequential)
always @(posedge clk) begin
    if(reg_write && rd != 0)
        regs[rd] <= wd;
end

endmodule
